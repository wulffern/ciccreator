*Testbench for SAR top level
*----------------------------------------------------------------------------
* OPTIONS
*----------------------------------------------------------------------------
.option method=gear gmin=1e-12 reltol=1e-6

*----------------------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------------------

.param vdd=1.6
.param vcm = 0.4

.param input_freq = 1e6

.param sample_width=25n
.param sample_period=100n
.param risefall = 1n
*----------------------------------------------------------------------------
* INCLUDES
*----------------------------------------------------------------------------
.include ../lay/SAR_ESSCIRC16_28N.spice
.include aimspice_model.spi

*----------------------------------------------------------------------------
* FORCE
*----------------------------------------------------------------------------
VDD AVDD 0 dc vdd
VSS AVSS 0 dc 0

VIP SAR_IP VCM SIN(0 0.4 input_freq 0 0) dc 0
VIN SAR_IN VCM SIN(0 -0.4 input_freq 0 0) dc 0
VCM VCM 0 dc vcm
VCK CK_SAMPLE 0 pulse(0 vdd 0 risefall risefall sample_width sample_period) dc 0

*----------------------------------------------------------------------------
* DUT
*----------------------------------------------------------------------------
XIV CK_SAMPLE EN AVDD AVSS IVX1_EV
XDUT SAR_IP SAR_IN SARN SARP DONE D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> EN CK_SAMPLE CK_SAMPLE AVDD AVDD AVSS SAR9B_EV


*----------------------------------------------------------------------------
* ANALYSIS
*----------------------------------------------------------------------------
.tran 1n 400n



