**********************************************************************
**        Copyright (c) 2014 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2014-5-9
** Author        : carsten (at) wulff.no
** *******************************************************************
**   Non-commercial use only, for commercial use contact license holder
**********************************************************************
**   This program is free software: you can redistribute it and/or modify
**   it under the terms of the GNU General Public License as published by
**   the Free Software Foundation, either version 3 of the License, or
**   (at your option) any later version.
** 
**   This program is distributed in the hope that it will be useful,
**   but WITHOUT ANY WARRANTY; without even the implied warranty of
**   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
**   GNU General Public License for more details.
** 
**   You should have received a copy of the GNU General Public License
**   along with this program.  If not, see <http://www.gnu.org/licenses/>.
**********************************************************************




*-----------------------------------------------------------------------------
* SAR unit logic cells
*---------------------------------------------------------------------------


.subckt TIEH_EV Y AVDD AVSS
MN0 A A AVSS AVSS NCHDL
MP0 Y A AVDD AVSS PCHDL
.ends TIEH_EV

.subckt TIEL_EV Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 A A AVDD AVSS PCHDL
.ends TIEL_EV

.subckt CAPX1_EV A B
XA1 A B CAPR
XB1 A B CAP
.ends

.subckt IVX1_EV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MP0 Y A AVDD AVSS PCHDL
.ends IVX1_EV

.subckt IVX2_EV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A AVDD AVSS PCHDL
MP1 AVDD A Y AVSS PCHDL
.ends IVX2_EV

.subckt IVX4_EV A Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A AVDD AVSS PCHDL
MP1 AVDD A Y AVSS PCHDL
MP2 Y A AVDD AVSS PCHDL
MP3 AVDD A Y AVSS PCHDL
.ends IVX4_EV

.subckt SWX2_EV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
.ends SWX2_EV

.SUBCKT TAPCELL_EV TAP
MN1 TAP TAP TAP TAP  NCHDL
MP1 TAP TAP TAP TAP  PCHDL
.ENDS

.subckt SWX4_EV A Y VREF AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS A Y AVSS NCHDL
MN2 Y A AVSS AVSS NCHDL
MN3 AVSS A Y AVSS NCHDL
MP0 Y A VREF AVSS PCHDL
MP1 VREF A Y AVSS PCHDL
MP2 Y A VREF AVSS PCHDL
MP3 VREF A Y AVSS PCHDL
.ends IVX4_EV

.subckt NRX1_EV A B Y AVDD AVSS
MN0 Y A AVSS AVSS NCHDL
MN1 AVSS B Y AVSS NCHDL
MP0 N1 A AVDD AVSS PCHDL
MP1 Y B N1 AVSS PCHDL
.ends NRX1_EV


.subckt NDX1_EV A B Y AVDD AVSS
MN0 N1 A AVSS AVSS NCHDL
MN1 Y B N1 AVSS NCHDL
MP0 Y A AVDD AVSS PCHDL
MP1 AVDD B Y AVSS PCHDL
.ends NDX1_EV

.subckt TGPD_EV C A B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN1 B C AVSS AVSS NCHDL
MN2 A CN B AVSS NCHDL
MP0 AVDD C CN AVSS PCHDL
MP1_DMY B AVDD AVDD AVSS PCHDL
MP2 A C B AVSS PCHDL
.ends

.subckt TAPCELLB_EV AVSS AVDD
MN1 AVSS AVSS AVSS AVSS  NCHDL
MP1 AVDD AVDD AVDD AVDD  PCHDL
.ends

.subckt SARBSSWCTRL_EV C GN GNG TIE_H  AVDD AVSS
MN0 N1 C AVSS AVSS NCHDL
MN1 GN TIE_H N1 AVSS NCHDL
MP0 GNG C GN AVSS PCHDL
MP1 AVDD GN GNG AVSS PCHDL
.ends

.SUBCKT SAREMX1_EV A  B EN ENO RST_N AVDD AVSS
MN0 N3 EN AM AVSS  NCHDL
MN1 N3 B AVSS AVSS  NCHDL
MN2 AVSS A N3 AVSS  NCHDL
MN3 ENO AM AVSS AVSS  NCHDL
MP0 AVDD RST_N AM AVSS PCHDL
MP1 N2 B ENO AVSS  PCHDL
MP2 N1 A N2 AVSS  PCHDL
MP3 AVDD AM N1 AVSS  PCHDL
.ENDS

.SUBCKT SARLTX1_EV A CHL RST_N EN LCK_N AVDD AVSS
MN0 N1 A AVSS AVSS  NCHDL
MN1 N3 LCK_N N1 AVSS  NCHDL
MN2 CHL EN N3 AVSS  NCHDL
MP0 NP2 RST_N AVDD AVSS PCHDL
MP1 NP1 RST_N NP2 AVSS PCHDL
MP2 CHL RST_N NP1 AVSS PCHDL
.ENDS

.SUBCKT SARCEX1_EV A B Y RST AVDD AVSS
MN0 N4 RST AVSS AVSS  NCHDL
MN1 AVSS RST N4 AVSS  NCHDL
MN2 N1 RST AVSS AVSS  NCHDL
MN3 Y RST N1 AVSS  NCHDL

MP0 N2 A Y AVSS PCHDL
MP1 AVDD A N2 AVSS PCHDL
MP2 N3 B AVDD AVSS PCHDL
MP3 Y B N3 AVSS PCHDL
.ENDS

.SUBCKT SARCMPHX1_EV CI CK CO VMR N1 N2 AVDD AVSS
MN0  N1 CK AVSS AVSS NCHDL
MN1  N2 CI N1   AVSS NCHDL
MN2  N1 CI N2   AVSS NCHDL
MN3  N2 CI N1   AVSS NCHDL
MN4  N1 CI N2   AVSS NCHDL
MN5  N2 CI N1   AVSS NCHDL
MN6  CO VMR N2   AVSS NCHDL

MP0  AVDD CK N1 AVSS PCHDL
MP1  N2 CK AVDD AVSS PCHDL
MP2  AVDD AVDD N2 AVSS PCHDL
MP3  CO CK AVDD AVSS PCHDL
MP4  AVDD VMR CO AVSS PCHDL
MP5  CO VMR AVDD AVSS PCHDL
MP6  AVDD VMR CO AVSS PCHDL
.ENDS SARCMPHX1_EV


.SUBCKT SARCMPHX2_EV CI CIR CK CO VMR N1 N2 AVDD AVSS
MN0  N1 CK AVSS AVSS NCHDL
MN1  N2 CI N1   AVSS NCHDL
MN2  N1 CI N2   AVSS NCHDL
MN3  N2 CI N1   AVSS NCHDL
MN4  N1 CI N2   AVSS NCHDL
MN3a  N2 CIR N1   AVSS NCHDL
MN4a  N1 CIR N2   AVSS NCHDL
MN3b  N2 CIR N1   AVSS NCHDL
MN4b  N1 CIR N2   AVSS NCHDL
MN5  N2 CIR N1   AVSS NCHDL
MN6  CO VMR N2   AVSS NCHDL

MP0  AVDD CK N1 AVSS PCHDL
MP1  N2 CK AVDD AVSS PCHDL
MP2  AVDD AVDD N2 AVSS PCHDL
MP2a  AVDD AVDD AVDD AVSS PCHDL
MP2b  AVDD AVDD AVDD AVSS PCHDL
MP2c  AVDD AVDD AVDD AVSS PCHDL
MP2d  AVDD AVDD AVDD AVSS PCHDL
MP3  CO CK AVDD AVSS PCHDL
MP4  AVDD VMR CO AVSS PCHDL
MP5  CO VMR AVDD AVSS PCHDL
MP6  AVDD VMR CO AVSS PCHDL

.ENDS SARCMPHX1_EV

.SUBCKT SARKICKHX1_EV CI CK CKN AVDD AVSS
MN0  N1 CKN AVSS AVSS NCHDL
MN1  N1 CI N1   AVSS NCHDL
MN2  N1 CI N1   AVSS NCHDL
MN3  N1 CI N1   AVSS NCHDL
MN4  N1 CI N1   AVSS NCHDL
MN5  N1 CI N1   AVSS NCHDL
MN6  AVDD CK N1   AVSS NCHDL

MP0  AVDD CKN N1 AVSS PCHDL
MP1_DMY AVDD AVDD AVDD AVSS PCHDL
MP2_DMY AVDD AVDD AVDD AVSS PCHDL
MP3_DMY AVDD AVDD AVDD AVSS PCHDL
MP4_DMY AVDD AVDD AVDD AVSS PCHDL
MP5_DMY AVDD AVDD AVDD AVSS PCHDL
MP6  AVDD AVDD AVDD AVSS PCHDL
.ENDS SARKICKHX1_EV

.SUBCKT SARKICKHX2_EV CI CIR CK CKN AVDD AVSS
MN0  N1 CKN AVSS AVSS NCHDL
MN1  N1 CI N1   AVSS NCHDL
MN2  N1 CI N1   AVSS NCHDL
MN3  N1 CI N1   AVSS NCHDL
MN4  N1 CI N1   AVSS NCHDL
MN3a  N1 CIR N1   AVSS NCHDL
MN4a  N1 CIR N1   AVSS NCHDL
MN3b  N1 CIR N1   AVSS NCHDL
MN4b  N1 CIR N1   AVSS NCHDL
MN5  N1 CIR N1   AVSS NCHDL
MN6  AVDD CK N1   AVSS NCHDL

MP0  AVDD CKN N1 AVSS PCHDL
MP1  AVDD AVDD AVDD AVSS PCHDL
MP2  AVDD AVDD AVDD AVSS PCHDL
MP3  AVDD AVDD AVDD AVSS PCHDL
MP4  AVDD AVDD AVDD AVSS PCHDL
MP3a  AVDD AVDD AVDD AVSS PCHDL
MP4a  AVDD AVDD AVDD AVSS PCHDL
MP3b  AVDD AVDD AVDD AVSS PCHDL
MP4b  AVDD AVDD AVDD AVSS PCHDL
MP5  AVDD AVDD AVDD AVSS PCHDL
MP6  AVDD AVDD AVDD AVSS PCHDL
.ENDS SARKICKHX2_EV


*-----------------------------------------------------------------------------
* SAR composite logic cells
*---------------------------------------------------------------------------


.SUBCKT SARBSSW_EV VI CK CKN TIE_L VO1 VO2 AVDD AVSS
M1 VI GN VO1 AVSS NCHDLR
M2 VI GN VO1 AVSS NCHDLR
M3 VI GN VO1 AVSS NCHDLR
M4 VI GN VO1 AVSS NCHDLR
M5 VI TIE_L VO2 AVSS NCHDLR
M6 VI TIE_L VO2 AVSS NCHDLR
M7 VI TIE_L VO2 AVSS NCHDLR
M8 VI TIE_L VO2 AVSS NCHDLR

XA0 CK CKN AVDD AVSS IVX1_EV
XA3 CKN VI VS AVDD AVSS TGPD_EV
XA4 CKN GN GNG TIE_H AVDD AVSS SARBSSWCTRL_EV
XA1 TIE_H AVDD AVSS TIEH_EV
XA2 TIE_L AVDD AVSS TIEL_EV
XA5 AVSS TAPCELL_EV
XCAPB GNG VS CAPX1_EV M=7
XCAPC GNG VS CAPX1_EV M=7

.ENDS

.SUBCKT SARCMPX1_EV CPI CNI CPO CNO CK_CMP CK_SAMPLE DONE AVDD AVSS
XA0 AVSS TAPCELL_EV
XA1 CPI CK_B CK_N AVDD AVSS SARKICKHX1_EV
XA2 CPI CK_B CNO_I CPO_I N1 NC1 AVDD AVSS SARCMPHX1_EV
XA2a CPO_I CPO AVDD AVSS IVX4_EV
XA3a CNO_I CNO AVDD AVSS IVX4_EV
XA3 CNI CK_B CPO_I CNO_I N1 NC2 AVDD AVSS SARCMPHX1_EV
XA4 CNI CK_B CK_N AVDD AVSS SARKICKHX1_EV
XA9 CK_N CK_B AVDD AVSS IVX1_EV
XA10 DONE_N CK_A CK_N AVDD AVSS NDX1_EV
XA11 CK_SAMPLE DONE DONE_N AVDD AVSS NRX1_EV
XA12 CK_CMP CK_A AVDD AVSS IVX1_EV
XA13 AVSS TAPCELL_EV
.ENDS


.SUBCKT SARMRYX1_EV CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS
XA0 AVSS TAPCELL_EV
XA1 CMP_OP CMP_ON EN ENO RST_N AVDD AVSS SAREMX1_EV
XA2 ENO LCK_N AVDD AVSS IVX1_EV
XA4 CMP_OP CHL_OP RST_N EN LCK_N AVDD AVSS SARLTX1_EV
XA5 CMP_ON CHL_ON RST_N EN LCK_N AVDD AVSS SARLTX1_EV
.ENDS

.SUBCKT SARDIGX1_EV CMP_OP CMP_ON EN RST_N ENO CP0 CP1 CN0 CN1 VREF AVDD AVSS
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON AVDD AVSS SARMRYX1_EV
XA2 CHL_ON CN1 VREF AVSS SWX2_EV
XA3 CN1 CP1 VREF AVSS SWX2_EV
XA4 CHL_OP CP0 VREF AVSS SWX2_EV
XA5 CP0 CN0 VREF AVSS SWX2_EV
XA6 AVSS TAPCELL_EV
.ENDS

.SUBCKT SARDIGEX2_EV CMP_OP CMP_ON EN RST_N ENO DONE CP0 CP1 CN0 CN1 CEIN CEO CKS VREF AVDD AVSS
XA1 CMP_OP CMP_ON EN RST_N ENO CHL_OP CHL_ON  AVDD AVSS SARMRYX1_EV

XA2 CHL_ON CN1 VREF AVSS SWX2_EV
XA3 CN1 CP1 VREF AVSS SWX2_EV
XA4 CHL_OP CP0 VREF AVSS SWX2_EV
XA5 CP0 CN0 VREF AVSS SWX2_EV

XA6 CN0 CP1 CE CKS AVDD AVSS SARCEX1_EV
XA7 ENO ENO_N AVDD AVSS IVX1_EV
XA8 ENO_N DONE AVDD AVSS IVX1_EV
XA9 ENO_N CE CE1 AVDD AVSS NDX1_EV
XA10 CE1 CE1_N AVDD AVSS IVX1_EV
XA11 CE1_N CEIN CEO1 AVDD AVSS NRX1_EV
XA12 CEO1 CEO AVDD AVSS IVX1_EV
XA13 AVSS TAPCELL_EV
.ENDS

*-----------------------------------------------------------------------------
* SAR capacitors
*-----------------------------------------------------------------------------


.subckt CAP32C_EV C1A C1B C2 C4 C8 C16 CTOP AVSS
*XR1 CTOP NCa RM4
*XR2 AVSS Ncb RM4

XRES1A C1A NC1 RM1
XRES1B C1B NC2 RM1
XRES2 C2 NC3 RM1
XRES4 C4 NC4 RM1
XRES8 C8 NC5 RM1
XRES16 C16 NC6 RM1
.ends CAP32C_EV


*-----------------------------------------------------------------------------
* SAR CDACs
*-----------------------------------------------------------------------------

.SUBCKT CDAC9_EV  CP<13> CP<12> CP<11> CP<10> CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0> CTOP  AVSS
XC1  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CAP32C_EV
XC256a<7>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CAP32C_EV
XC128b<3>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CAP32C_EV
XC64a<0>  CP<8> CP<8> CP<8> CP<8> CP<8> CP<8> CTOP AVSS  CAP32C_EV
XC32a<0>  CP<6> CP<6> CP<6> CP<6> CP<6> CP<7> CTOP AVSS  CAP32C_EV
XCS       AVSS CP<0> CP<1> CP<2> CP<3>  AVSS CTOP AVSS  CAP32C_EV
XC128a<1>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CAP32C_EV
XC256b<5>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CAP32C_EV
XC256a<5>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CAP32C_EV
XC256b<2>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CAP32C_EV
XC256a<2>  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CAP32C_EV
XC128b<2>  CP<10> CP<10> CP<10> CP<10> CP<10> CP<10> CTOP AVSS  CAP32C_EV
X16ab       CP<5> CP<5> CP<5> CP<5> CP<4> AVSS CTOP AVSS  CAP32C_EV
XC64b<1>  CP<9> CP<9> CP<9> CP<9> CP<9> CP<9> CTOP AVSS  CAP32C_EV
XC128a<0>  CP<11> CP<11> CP<11> CP<11> CP<11> CP<11> CTOP AVSS  CAP32C_EV
XC256b<0>  CP<12> CP<12> CP<12> CP<12> CP<12> CP<12> CTOP AVSS  CAP32C_EV
XC0  CP<13> CP<13> CP<13> CP<13> CP<13> CP<13> CTOP AVSS  CAP32C_EV
.ENDS CDAC9_EV

*-----------------------------------------------------------------------------
* SAR CDACs with logic
*-----------------------------------------------------------------------------

.SUBCKT SAR9B_EV_NOROUTE SAR_IP SAR_IN SARN SARP DONE D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> EN CK_SAMPLE  CK_SAMPLE_BSSW  VREF AVDD AVSS

XB1  SAR_IP CK_SAMPLE_BSSW NCCA CEIN SARP SARN AVDD AVSS SARBSSW_EV
XB2  SAR_IN CK_SAMPLE_BSSW NCCB CEIN SARN SARP AVDD AVSS SARBSSW_EV

XDAC1  CP<13> CP<12> D<8> CP<10> D<7> CP<8> D<6> CP<6> D<5> CP<4> D<4> D<3> D<2> D<1> SARP AVSS CDAC9_EV
XDAC2  D<9> CN<12> CN<11> CN<10> CN<9> CN<8> CN<7> CN<6> CN<5> CN<4> CN<3> CN<2> CN<1> CN<0> SARN  AVSS CDAC9_EV

XA0 CMP_OP CMP_ON EN EN ENO0 DONE0 CP<12> CP<13> CN<12> D<9> CEIN CEO0 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA1 CMP_OP CMP_ON ENO0 EN ENO1 DONE1 CP<10> D<8> CN<10> CN<11> CEO0 CEO1 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA2 CMP_OP CMP_ON ENO1 EN ENO2 DONE2 CP<8> D<7> CN<8> CN<9> CEO1 CEO2 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA3 CMP_OP CMP_ON ENO2 EN ENO3 DONE3 CP<6> D<6> CN<6> CN<7> CEO2 CEO3 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA4 CMP_OP CMP_ON ENO3 EN ENO4 DONE4 CP<4> D<5> CN<4> CN<5> CEO3 CEO4 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA5 CMP_OP CMP_ON ENO4 EN ENO5 DONE5 NC3A D<4> CN<3> NC3B CEO4 CEO5 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA6 CMP_OP CMP_ON ENO5 EN ENO6 DONE6 NC4A D<3> CN<2> NC4B CEO5 CEO6 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA7 CMP_OP CMP_ON ENO6 EN ENO7 DONE7 NC5A D<2> CN<1> NC5B CEO6 CEO7 CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV
XA8 CMP_OP CMP_ON ENO7 EN ENO8 DONE NC6A D<1> CN<0> NC6B CEO7 CK_CMP CK_SAMPLE VREF AVDD AVSS SARDIGEX4_EV

XA20 SARP SARN CMP_OP CMP_ON CK_CMP CK_SAMPLE DONE AVDD AVSS SARCMPX1_EV
.ENDS
