*Test model for use with eldo and cIcCreator
.model nch NMOS level=60
.model nch_lvt NMOS level=60
.model nch_io NMOS level=60
.model nch_lvt_io NMOS level=60

.model pch PMOS level=60 
.model pch_lvt PMOS level=60
.model pch_io PMOS level=60
.model pch_lvt_io PMOS level=60


