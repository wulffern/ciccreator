*Testbench for boostrapped switch
*----------------------------------------------------------------------------
* OPTIONS
*----------------------------------------------------------------------------
.option method=gear gmin=1e-12 reltol=1e-6

*----------------------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------------------

.param vdd=1.6
.param vcm = 0.4

.param input_freq = 1e5

.param cmp_width=200n
.param cmp_period=400n
.param risefall = 1n
*----------------------------------------------------------------------------
* INCLUDES
*----------------------------------------------------------------------------
.include ../lay/SAR_ESSCIRC16_28N.spice
.include aimspice_model.spi

*----------------------------------------------------------------------------
* FORCE
*----------------------------------------------------------------------------
VDD AVDD 0 dc vdd
VSS AVSS 0 dc 0

VIP SAR_IP VCM SIN(0 0.4 input_freq 0 0) dc 0
VIN SAR_IN VCM SIN(0 -0.4 input_freq 0 0) dc 0
VCM VCM 0 dc vcm
VCK CK_SAMPLE 0 dc 0
VDONE DONE 0 dc 0
VCMP CK_CMP 0 pulse(0 vdd 0 risefall risefall cmp_width cmp_period) dc 0

*----------------------------------------------------------------------------
* DUT
*----------------------------------------------------------------------------
XA20 SAR_IP SAR_IN CMP_OP CMP_ON CK_CMP CK_SAMPLE DONE AVDD AVSS SARCMPX1_EV 




*----------------------------------------------------------------------------
* ANALYSIS
*----------------------------------------------------------------------------
.tran 1n 10u



