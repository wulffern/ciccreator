*Testbench for boostrapped switch
*----------------------------------------------------------------------------
* OPTIONS
*----------------------------------------------------------------------------
.option method=gear gmin=1e-12 reltol=1e-6


*----------------------------------------------------------------------------
* PARAMETERS
*----------------------------------------------------------------------------

.param vdd=1.6
.param vcm = 0.4

.param input_freq = 1e6

.param sample_width=10n
.param sample_period=40n
.param risefall = 1n

*----------------------------------------------------------------------------
* INCULDE
*----------------------------------------------------------------------------
.include model.spi


*----------------------------------------------------------------------------
* DUT
*----------------------------------------------------------------------------
XB1 SAR_IP CK_SAMPLE NCCA CEIN SARP SARN AVDD AVSS SARBSSW_EV
XB2 SAR_IN CK_SAMPLE NCCB CEIN SARN SARP AVDD AVSS SARBSSW_EV 

C1 SARP 0 0.5p
C2 SARN 0 0.5p



*----------------------------------------------------------------------------
* FORCE
*----------------------------------------------------------------------------
VDD AVDD 0 dc vdd
VSS AVSS 0 dc 0

VIP SAR_IP VCM SIN(0 0.4 input_freq 0 0) dc 0
VIN SAR_IN VCM SIN(0 -0.4 input_freq 0 0) dc 0
VCM VCM 0 dc vcm
VCK CK_SAMPLE 0 pulse(0 vdd 0 risefall risefall sample_width sample_period) dc 0

bin vi 0 v=(v(SAR_IP) - v(SAR_IN))
bon vo 0 v=(v(sarp) - v(sarn))
*----------------------------------------------------------------------------
* ANALYSIS
*----------------------------------------------------------------------------
.tran 1n 2u

*----------------------------------------------------------------------------
* PLOTS AND EXTRACTS
*----------------------------------------------------------------------------
.plot v(SAR_IP) v(SARP) v(SAR_IN) v(SARN)
.plot v(CK_SAMPLE)
.plot v(vi) v(vo)

